library verilog;
use verilog.vl_types.all;
entity ins_ram_tb is
end ins_ram_tb;
