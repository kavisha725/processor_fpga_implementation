library verilog;
use verilog.vl_types.all;
entity img_in_ddr_tb is
end img_in_ddr_tb;
